module team_06_reverb (
    input logic clk, rst,
    input logic audio_in,
    output logic reverb_out
);




endmodule