module i2sclock (
    input logic clk, rst,
    output curr_i2sclk, past_i2sclk
);
endmodule