module display
( 
    input logic state,
    output logic lcdData
);



endmodule;