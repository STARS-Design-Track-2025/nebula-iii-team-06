module team_06_edge_detection_i2s(
    input logic i2sclk,
    output logic curr_i2sclk, past_i2sclk
);
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            curr_i2sclk <= 0;
            past_i2sclk <= 0;
        end else begin
            past_i2sclk <= curr_i2sclk;
            curr_i2sclk <= i2s_sck;
        end
end
endmodule